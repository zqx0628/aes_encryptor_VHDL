library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package util_package is    
    function mtp2 (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function mtpe (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function mtpb (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function mtpd (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function mtp9 (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function sbox (x:std_logic_vector(7 downto 0)) return std_logic_vector;
    function T (j:integer;x:std_logic_vector(31 downto 0)) return std_logic_vector;
end util_package;

package body util_package is

function mtp2 (x : std_logic_vector(7 downto 0)) return std_logic_vector is
    variable i : std_logic_vector(7 downto 0);
begin
    if x(7)='0' then
        i:=x(6 downto 0)&"0";
    else
        i:=(x(6 downto 0)&"0") xor "00011011";
    end if;
    return i;
end function;

function mtpe (x:std_logic_vector(7 downto 0)) return std_logic_vector is
begin
    return mtp2(mtp2(mtp2(x))) xor mtp2(mtp2(x)) xor mtp2(x);
end function;

function mtpb (x:std_logic_vector(7 downto 0)) return std_logic_vector is
begin
    return mtp2(mtp2(mtp2(x))) xor mtp2(x) xor x;
end function;

function mtpd (x:std_logic_vector(7 downto 0)) return std_logic_vector is
begin
    return mtp2(mtp2(mtp2(x))) xor mtp2(mtp2(x)) xor x;
end function;

function mtp9 (x:std_logic_vector(7 downto 0)) return std_logic_vector is
begin
    return mtp2(mtp2(mtp2(x))) xor x;
end function;

function T (j:integer;x:std_logic_vector(31 downto 0)) return std_logic_vector is
    variable a:std_logic_vector(31 downto 0);
    variable b:std_logic_vector(31 downto 0);
    variable c:std_logic_vector(31 downto 0);
begin
    a:=x(23 downto 0)&x(31 downto 24);
    b:=sbox(a(31 downto 24)) & sbox(a(23 downto 16)) & sbox(a(15 downto 8)) & sbox(a(7 downto 0));
    case j is
        when 1 => c:= "00000001000000000000000000000000" xor b;
        when 2 => c:= "00000010000000000000000000000000" xor b;
        when 3 => c:= "00000100000000000000000000000000" xor b;
        when 4 => c:= "00001000000000000000000000000000" xor b;
        when 5 => c:= "00010000000000000000000000000000" xor b;
        when 6 => c:= "00100000000000000000000000000000" xor b;
        when 7 => c:= "01000000000000000000000000000000" xor b;
        when 8 => c:= "10000000000000000000000000000000" xor b;
        when 9 => c:= "00011011000000000000000000000000" xor b;
        when 10=> c:= "00110110000000000000000000000000" xor b;
        when others => c:="00000000000000000000000000000000";
    end case;
    return c;
end function;

function sbox (x: std_logic_vector(7 downto 0)) return std_logic_vector is 
    variable i:std_logic_vector(7 downto 0);
begin
    case x is
        when "00000000" =>i:="01100011";
		when "00000001" =>i:="01111100";
		when "00000010" =>i:="01110111";
		when "00000011" =>i:="01111011";
		when "00000100" =>i:="11110010";
		when "00000101" =>i:="01101011";
		when "00000110" =>i:="01101111";
		when "00000111" =>i:="11000101";
		when "00001000" =>i:="00110000";
		when "00001001" =>i:="00000001";
		when "00001010" =>i:="01100111";
		when "00001011" =>i:="00101011";
		when "00001100" =>i:="11111110";
		when "00001101" =>i:="11010111";
		when "00001110" =>i:="10101011";
		when "00001111" =>i:="01110110";
		when "00010000" =>i:="11001010";
		when "00010001" =>i:="10000010";
		when "00010010" =>i:="11001001";
		when "00010011" =>i:="01111101";
		when "00010100" =>i:="11111010";
		when "00010101" =>i:="01011001";
		when "00010110" =>i:="01000111";
		when "00010111" =>i:="11110000";
		when "00011000" =>i:="10101101";
		when "00011001" =>i:="11010100";
		when "00011010" =>i:="10100010";
		when "00011011" =>i:="10101111";
		when "00011100" =>i:="10011100";
		when "00011101" =>i:="10100100";
		when "00011110" =>i:="01110010";
		when "00011111" =>i:="11000000";
		when "00100000" =>i:="10110111";
		when "00100001" =>i:="11111101";
		when "00100010" =>i:="10010011";
		when "00100011" =>i:="00100110";
		when "00100100" =>i:="00110110";
		when "00100101" =>i:="00111111";
		when "00100110" =>i:="11110111";
		when "00100111" =>i:="11001100";
		when "00101000" =>i:="00110100";
		when "00101001" =>i:="10100101";
		when "00101010" =>i:="11100101";
		when "00101011" =>i:="11110001";
		when "00101100" =>i:="01110001";
		when "00101101" =>i:="11011000";
		when "00101110" =>i:="00110001";
		when "00101111" =>i:="00010101";
		when "00110000" =>i:="00000100";
		when "00110001" =>i:="11000111";
		when "00110010" =>i:="00100011";
		when "00110011" =>i:="11000011";
		when "00110100" =>i:="00011000";
		when "00110101" =>i:="10010110";
		when "00110110" =>i:="00000101";
		when "00110111" =>i:="10011010";
		when "00111000" =>i:="00000111";
		when "00111001" =>i:="00010010";
		when "00111010" =>i:="10000000";
		when "00111011" =>i:="11100010";
		when "00111100" =>i:="11101011";
		when "00111101" =>i:="00100111";
		when "00111110" =>i:="10110010";
		when "00111111" =>i:="01110101";
		when "01000000" =>i:="00001001";
		when "01000001" =>i:="10000011";
		when "01000010" =>i:="00101100";
		when "01000011" =>i:="00011010";
		when "01000100" =>i:="00011011";
		when "01000101" =>i:="01101110";
		when "01000110" =>i:="01011010";
		when "01000111" =>i:="10100000";
		when "01001000" =>i:="01010010";
		when "01001001" =>i:="00111011";
		when "01001010" =>i:="11010110";
		when "01001011" =>i:="10110011";
		when "01001100" =>i:="00101001";
		when "01001101" =>i:="11100011";
		when "01001110" =>i:="00101111";
		when "01001111" =>i:="10000100";
		when "01010000" =>i:="01010011";
		when "01010001" =>i:="11010001";
		when "01010010" =>i:="00000000";
		when "01010011" =>i:="11101101";
		when "01010100" =>i:="00100000";
		when "01010101" =>i:="11111100";
		when "01010110" =>i:="10110001";
		when "01010111" =>i:="01011011";
		when "01011000" =>i:="01101010";
		when "01011001" =>i:="11001011";
		when "01011010" =>i:="10111110";
		when "01011011" =>i:="00111001";
		when "01011100" =>i:="01001010";
		when "01011101" =>i:="01001100";
		when "01011110" =>i:="01011000";
		when "01011111" =>i:="11001111";
		when "01100000" =>i:="11010000";
		when "01100001" =>i:="11101111";
		when "01100010" =>i:="10101010";
		when "01100011" =>i:="11111011";
		when "01100100" =>i:="01000011";
		when "01100101" =>i:="01001101";
		when "01100110" =>i:="00110011";
		when "01100111" =>i:="10000101";
		when "01101000" =>i:="01000101";
		when "01101001" =>i:="11111001";
		when "01101010" =>i:="00000010";
		when "01101011" =>i:="01111111";
		when "01101100" =>i:="01010000";
		when "01101101" =>i:="00111100";
		when "01101110" =>i:="10011111";
		when "01101111" =>i:="10101000";
		when "01110000" =>i:="01010001";
		when "01110001" =>i:="10100011";
		when "01110010" =>i:="01000000";
		when "01110011" =>i:="10001111";
		when "01110100" =>i:="10010010";
		when "01110101" =>i:="10011101";
		when "01110110" =>i:="00111000";
		when "01110111" =>i:="11110101";
		when "01111000" =>i:="10111100";
		when "01111001" =>i:="10110110";
		when "01111010" =>i:="11011010";
		when "01111011" =>i:="00100001";
		when "01111100" =>i:="00010000";
		when "01111101" =>i:="11111111";
		when "01111110" =>i:="11110011";
		when "01111111" =>i:="11010010";
		when "10000000" =>i:="11001101";
		when "10000001" =>i:="00001100";
		when "10000010" =>i:="00010011";
		when "10000011" =>i:="11101100";
		when "10000100" =>i:="01011111";
		when "10000101" =>i:="10010111";
		when "10000110" =>i:="01000100";
		when "10000111" =>i:="00010111";
		when "10001000" =>i:="11000100";
		when "10001001" =>i:="10100111";
		when "10001010" =>i:="01111110";
		when "10001011" =>i:="00111101";
		when "10001100" =>i:="01100100";
		when "10001101" =>i:="01011101";
		when "10001110" =>i:="00011001";
		when "10001111" =>i:="01110011";
		when "10010000" =>i:="01100000";
		when "10010001" =>i:="10000001";
		when "10010010" =>i:="01001111";
		when "10010011" =>i:="11011100";
		when "10010100" =>i:="00100010";
		when "10010101" =>i:="00101010";
		when "10010110" =>i:="10010000";
		when "10010111" =>i:="10001000";
		when "10011000" =>i:="01000110";
		when "10011001" =>i:="11101110";
		when "10011010" =>i:="10111000";
		when "10011011" =>i:="00010100";
		when "10011100" =>i:="11011110";
		when "10011101" =>i:="01011110";
		when "10011110" =>i:="00001011";
		when "10011111" =>i:="11011011";
		when "10100000" =>i:="11100000";
		when "10100001" =>i:="00110010";
		when "10100010" =>i:="00111010";
		when "10100011" =>i:="00001010";
		when "10100100" =>i:="01001001";
		when "10100101" =>i:="00000110";
		when "10100110" =>i:="00100100";
		when "10100111" =>i:="01011100";
		when "10101000" =>i:="11000010";
		when "10101001" =>i:="11010011";
		when "10101010" =>i:="10101100";
		when "10101011" =>i:="01100010";
		when "10101100" =>i:="10010001";
		when "10101101" =>i:="10010101";
		when "10101110" =>i:="11100100";
		when "10101111" =>i:="01111001";
		when "10110000" =>i:="11100111";
		when "10110001" =>i:="11001000";
		when "10110010" =>i:="00110111";
		when "10110011" =>i:="01101101";
		when "10110100" =>i:="10001101";
		when "10110101" =>i:="11010101";
		when "10110110" =>i:="01001110";
		when "10110111" =>i:="10101001";
		when "10111000" =>i:="01101100";
		when "10111001" =>i:="01010110";
		when "10111010" =>i:="11110100";
		when "10111011" =>i:="11101010";
		when "10111100" =>i:="01100101";
		when "10111101" =>i:="01111010";
		when "10111110" =>i:="10101110";
		when "10111111" =>i:="00001000";
		when "11000000" =>i:="10111010";
		when "11000001" =>i:="01111000";
		when "11000010" =>i:="00100101";
		when "11000011" =>i:="00101110";
		when "11000100" =>i:="00011100";
		when "11000101" =>i:="10100110";
		when "11000110" =>i:="10110100";
		when "11000111" =>i:="11000110";
		when "11001000" =>i:="11101000";
		when "11001001" =>i:="11011101";
		when "11001010" =>i:="01110100";
		when "11001011" =>i:="00011111";
		when "11001100" =>i:="01001011";
		when "11001101" =>i:="10111101";
		when "11001110" =>i:="10001011";
		when "11001111" =>i:="10001010";
		when "11010000" =>i:="01110000";
		when "11010001" =>i:="00111110";
		when "11010010" =>i:="10110101";
		when "11010011" =>i:="01100110";
		when "11010100" =>i:="01001000";
		when "11010101" =>i:="00000011";
		when "11010110" =>i:="11110110";
		when "11010111" =>i:="00001110";
		when "11011000" =>i:="01100001";
		when "11011001" =>i:="00110101";
		when "11011010" =>i:="01010111";
		when "11011011" =>i:="10111001";
		when "11011100" =>i:="10000110";
		when "11011101" =>i:="11000001";
		when "11011110" =>i:="00011101";
		when "11011111" =>i:="10011110";
		when "11100000" =>i:="11100001";
		when "11100001" =>i:="11111000";
		when "11100010" =>i:="10011000";
		when "11100011" =>i:="00010001";
		when "11100100" =>i:="01101001";
		when "11100101" =>i:="11011001";
		when "11100110" =>i:="10001110";
		when "11100111" =>i:="10010100";
		when "11101000" =>i:="10011011";
		when "11101001" =>i:="00011110";
		when "11101010" =>i:="10000111";
		when "11101011" =>i:="11101001";
		when "11101100" =>i:="11001110";
		when "11101101" =>i:="01010101";
		when "11101110" =>i:="00101000";
		when "11101111" =>i:="11011111";
		when "11110000" =>i:="10001100";
		when "11110001" =>i:="10100001";
		when "11110010" =>i:="10001001";
		when "11110011" =>i:="00001101";
		when "11110100" =>i:="10111111";
		when "11110101" =>i:="11100110";
		when "11110110" =>i:="01000010";
		when "11110111" =>i:="01101000";
		when "11111000" =>i:="01000001";
		when "11111001" =>i:="10011001";
		when "11111010" =>i:="00101101";
		when "11111011" =>i:="00001111";
		when "11111100" =>i:="10110000";
		when "11111101" =>i:="01010100";
		when "11111110" =>i:="10111011";
		when "11111111" =>i:="00010110";
        when others=>i:="00000000";
    end case;
    return i;
end function;
end package body util_package;